interface tb_interface(input logic clk);
logic rst;
logic [63:0] rx_data_net;
logic [6:0] counterOut;
logic [47:0] dMac_out;
logic [47:0] sMac_out;
logic [15:0] oTag_out;
logic [15:0] eType_out;
logic [3:0] version_out;
logic [3:0] headerLength_out;
logic [7:0] typeOfService_out;
logic [15:0] totalLength_out;
logic [15:0] identification_out;
logic [2:0] flags_out;
logic [12:0] fragmentOffset_out;
logic [7:0] timeToLive_out;
logic [7:0] protocol_out;
logic [15:0] headerChecksum_out;
logic [31:0] srcIPAddress_out;
logic [31:0] destIPAddress_out;
logic [15:0] srcPort_out;
logic [15:0] destPort_out;
logic [15:0] length_out;
logic [15:0] checksum_out;
logic [79:0] sessionID_out;
logic [63:0] sequenceNumber_out;
logic [15:0] messageCount_out;
clocking cb @(posedge clk);
    default input #1step output#3;
    //output rst;
    output  rx_data_net;
    input  counterOut;
    input  dMac_out;
    input sMac_out;
    input oTag_out;
    input eType_out;
    input version_out;
    input headerLength_out;
    input typeOfService_out;
    input totalLength_out;
    input identification_out;
    input flags_out;
    input fragmentOffset_out;
    input timeToLive_out;
    input protocol_out;
    input headerChecksum_out;
    input srcIPAddress_out;
    input destIPAddress_out;
    input srcPort_out;
    input destPort_out;
    input length_out;
    input checksum_out;
    input sessionID_out;
    input sequenceNumber_out;
    input messageCount_out;
endclocking
endinterface //tb_interface